Här är Freetype Manager, som används för att installera och konfigurera
nya Truetype-typsnitt i systemet. Inte så användarvänligt, men du kan pilla
på varje liten detalj. Ännu viktigare, det fungerar. :-)
