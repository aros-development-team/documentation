.. raw:: html

   <div class="front-container">

   <div class="main-div"><!--left side with main content-->

   <section>

.. Include:: introduction/index-abstract.sv

`Läs mer... <introduction/index>`__

.. raw:: html

   </section>

   <section>

   <h1>Distributioner<br><img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"></h1>

.. Include:: download-abstract.sv

`Läs mer... <download>`__

.. raw:: html

   </section>

   <section>

   <h1>GitHub Commits<br><img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"></h1>
   <object width="100%" height="250" data="github-commits.php" type="text/html"></object>

   </section>

   <section>

.. Include:: news/index.sv

.. raw:: html

   </section>

   </div><!--main-div-->

   <div class="rss-div"><!--right side with rss feeds-->

   <div class="rssfeed">

   <img alt="Archive Icon" src="/images/archivedownloadicon.png" align="top"><br>
   Latest ARCHIVE submissions:<br>
   <img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"><br>
   På <a href=https://archives.arosworld.org>The AROS archives</a>
   hittar du det nyaste materialet för AROS, här hittar du program, teman, grafik och ytterligare dokumentation.<br><br>
   <object width="100%" height="300" data="archives-uploads.php" type="text/html"></object>

   </div>

   <div class="rssfeed">

   <img alt="Community Icon" src="/images/communityicon.png" align="top"><br>
   Senaste inläggen på AROSWorld forumet:<br>
   <img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"><br>
   <a href=https://www.arosworld.org>AROSWorld</a>
   är den primära AROS community-sidan. Här kan du få hjälp, hålla koll på vad som händer inom AROS-världen och posta dina tankar om AROS.<br><br>
   <object width="100%" height="400" data="arosworld-forum.php" type="text/html"></object>

   </div>

   </div><!--rss-div-->
   </div><!--front-container-->
