.. raw:: html

   <h1>Distributioner<br><img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"></h1>

Detta �r f�rkonfigurerade och v�ltestade versioner av AROS. De inneh�ller
m�nga anv�ndbara program som inte f�ljer med fr�n start och �r de som �r mest
intressanta f�r vanliga anv�ndare. De kanske saknar den senaste versionen av
AROS, men de �r mycket stabilare och mer anv�ndarv�nliga �n nightly builds.
Om du �r en som �r nyfiken p� vad AROS har att erbjuda s� rekommenderar vi att
du anv�nder distributioner f�r b�sta m�jliga upplevelse.

