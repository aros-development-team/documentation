Sponsorer
=========

:Authors:   Aaron Digulla, Adam Chodorowski 
:Copyright: Copyright © 1995-2002, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.


Följande företag, organisationer och individer har donerat resurser:

+ Trustec__
   
  .. RAW:: html
     
     <a href="http://www.trustsec.de/"><img border="0" src="/images/trustec.png"></a>
    
  De snälla personerna på Trustec donerar utrymme och bandbredd till AROS
  webbserver, SVN-server, FTP-server och flera mailinglistor. Om du är i behov
  av Java-utveckling eller kurser i Tyskland, kontakta dem!

+ Genesi__

  .. RAW:: html
  
     <a href="http://www.pegasosppc.com/"><img border="0" src="/images/genesi.gif"></a>

  Genesi har varit generösa och donerat ett Pegasos moderkort för att möjliggöra ett
  försök att porta AROS till den plattforman, tack!

+ SourceForge__

  .. RAW:: html
  
     <a href="http://www.sourceforge.net/"><img border="0" src="/images/sourceforge.png"></a>

  SourceForge försörjer oss med flera tjänster, såsom webbserver med möjligheter
  att köra skript, SQL-databas, mailinglistor, buggdatabas och ett distribuerat
  system för distribution av filer.

+ Yann Vernier
+ Randal Vice


Följande organisationer och individer har sponsrat utvecklingsarbete:

+ `Team AROS`__
+ `Norsk Amigaforening`__
+ Timothy Rue
+ Jakob Eriksson
+ Serge Guillaume
+ David Ferguson
+ Nils-Erik Reklev Skilnand
+ Jonny Johansson
+ Johan Grip
+ Marcus Karlsson
+ Rune Jensen
+ Joshua Dolan
+ Matthew Parsons
+ Jean-Pierre Rivière

__ http://www.trustsec.de/
__ http://www.pegasosppc.com/
__ http://www.sourceforge.net/
__ http://www.thenostromo.com/teamaros/
__ http://www.naf.as/
