.. raw:: html

   <h1>Introduktion<br><img style="width: 238px; height: 2px;" alt="" src="/images/sidespacer.png" /></h1>

.. raw:: html

  <?php include('/home/project-web/aros/htdocs/rsfeed/randimg.php');  random_image("/images/thubs/","100","76"); ?>

AROS �r ett resurssn�lt, effektivt och flexibelt operativsystem, gjord f�r att
hj�lpa dig f� ut det mesta av din dator. Det �r ett oberoende, fritt och
plattforms�verskridande projekt med m�let att vara kompatibelt med AmigaOS p�
API-niv� (p� samma s�tt som Wine, men olikt UAE), men f�rb�ttrat p� flertalet
omr�den. K�llkoden �r tillg�nglig under en "�ppen-k�llkod"-licens vilket
till�ter att vem som helst f�r g�ra f�rb�ttringar.

