Tids-inställnings-applikationen, klockan och WritePixelArrayAlpha testprogrammen
som visar alpha blending.
