========
Länkning
========

:Author:    Adam Chodorowski
:Copyright: Copyright Š 2001-2007, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.

Ett mycket bra sätt att visa ditt stöd för AROS, och för att uppmana andra,
är att länka till denna hemsida från din egen. Du kan använda en av nedanstående banners
för detta ändamål.

+------------------------------------------+----------------------+
| Bild                                     | Upphovsman           |
+==========================================+======================+
| .. Image:: /images/aros-banner.gif       | Cyb0rg / Resistance  |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner2.png      | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-blue.png  | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-pb2.png   | Paolo Besser         |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-banner-peta.png  | Petr Novak           |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+


Alternativt så finns det även signatur-banners för användning i forum:

+------------------------------------------+----------------------+
| Bild                                     | Upphovsman           |
+==========================================+======================+
| .. Image:: /images/aros-sigbar-user.png  | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+
| .. Image:: /images/aros-sigbar-coder.png | S33k_100             |
|  :align: center                          |                      |
|  :class: bannerimage                     |                      |
+------------------------------------------+----------------------+


Var vänlig, länka direkt till http://www.aros.org/ och inte till någon av de speglade
hemsidorna eftersom dessa kan ändras. Se även till att ha en lokal kopia av bilden för
att minska bandbredden.
