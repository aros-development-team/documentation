=============
Status Update
=============

:Author:   Paolo Besser
:Date:     2007-10-01

Senaste nyheter
---------------

Nyhet! Neil Cafferkey har bidragit med en helt ny `installer`__ för
AROS, vilket möjliggör en renare och säkrare installation på hårddiskar.
Nya finnesser enligt nedan:

- Installationsdisk och partitioner kan nu anges.
- Skapandet av en Work-partition fungerar.
- Partitionsstorlekar kan anges och existerande partitioner kan behållas.
- Windows är tillagd till GRUB boot menu om en existerande Windows-partition hittas.


Notera dock, att detta fortfarande är en beta-version. Här följer några
varningar från Neil: " Den nya hårddisk-installern är nu inkluderad
i "Nightly ISO" och är färdig för testning. Men, det finns för tillfället
en bug i antingen Wanderer eller FFS som måste åtgärdas. Efter att man startat
installern, så måste du avsluta Wanderer innan du fortsätter (om du inte
kommer att formatera någon partition).
Var extra försiktig än vanligt med denna version av installern, utsätt inte
datorn med ej säkerhetskopierad data. Den borde behålla alla existerande
partitioner, men inte så många har testat detta förutom jag."

Om du har en testdator med ej viktig data på, så vore det bästa om du
laddar ner 10-01 "nightly build (eller senare) och hjälper oss att hitta
buggar. Du kan använda Bug Tracker eller skicka ett meddelande i detta
AROS-Exec `discussion`__. 

Demonstration av AROS
---------------------

Som tidigare nämnt på denna hemsida så har AROS varit en gäststjärna på
`Pianeta Amiga 2007`__.  Under den populära amigashowen så har
Paulo Besser presenterat AROS till en del intresserade Amiga-anhängare.
Evenemanget har nämnts i några större IT-nyhets-hemsidor som `TGM Online`__
och `HW Upgrade`__. En rapport av evenemanget har blivit publicerad av 
`The AROS Show`__ (Läs denna `here`__) Du kan även se en trevlig `video`__
på YouTube.

__ http://mama.indstate.edu/users/nova/installer.jpg
__ https://ae.amigalife.org/modules/newbb/viewtopic.php?topic_id=2319
__ http://www.pianetaamiga.it/2007/eng/
__ http://tgmonline.futuregamer.it/news/settembre2007/20070910111905
__ http://www.hwupgrade.it/news/videogiochi/presentazione-italiana-per-l-os-indipendente-aros_22619-0.html
__ http://arosshow.blogspot.com
__ http://arosshow.blogspot.com/2007/09/pianeta-amiga-2007-report-from-paolo.html
__ http://video.google.it/videoplay?docid=-3563710058663289244
