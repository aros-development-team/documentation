Zune blir bara bättre och bättre! Nu tack vare Georg Steger så har
vi fler classes implementerade, som du kan se. Du kan även se gcc
kompilera ett av test-programmen för de nya implementerade classes.
