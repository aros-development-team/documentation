Mer sidor i Zune-inställningarna.
