.. raw:: html

   <h1>Distributioner<br><img style="width: 238px; height: 2px;" alt="spacer" src="/images/sidespacer.png"></h1>

Detta är förkonfigurerade och vältestade versioner av AROS. De innehåller
många användbara program som inte följer med från start och är de som är mest
intressanta för vanliga användare. De kanske saknar den senaste versionen av
AROS, men de är mycket stabilare och mer användarvänliga än nightly builds.
Om du är en som är nyfiken på vad AROS har att erbjuda så rekommenderar vi att
du använder distributioner för bästa möjliga upplevelse.

