Mer sidor i Zune-inställningar, så du kan konfigurera användarinterfacet
precis som *du* vill ha det.
