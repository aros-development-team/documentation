Här har vi några nya funktioner i icon-library. Du kan se den nya effekten 
för de valda ikonerna ("S"-mappen är vald här, därför är den ljusare än de
andra ikonerna). Ikon-namnen ritas nu upp med en outline, för att bli 
synliga även på en mörk bakgrund (detta kommer naturligtvis även att vara
konfigurerbart för användarna i framtiden).

Vi kan även se fil-identifikationen i bruk: text-filerna i "S"-mappen får
speciella def_Text-ikoner, medans filen "AROS.png" får den generella
projekt-ikonen. Vi har inte så många ikoner just nu, men om de fanns
tillgängliga så skulle "AROS.png" få en def_Picture-ikon (Eller även kanske
en def_PNG-ikon om det fanns tillgängligt).
