=================
Statusuppdatering
=================

:Författare:   Paolo Besser
:Datum:     2006-09-15

Översättningen av aros.org fortsätter. Samuel Atlan jobbar på sin
`Franska översättning`__ av vår hemsida. Det kommer att ta lite tid
innan det blir färdigt men de första sidorna finns redans tillgängliga
från menyn i övre vänstra hörnet. Nytt på aros.org är också att man
nu kan nå de översatta sidorna genom att lägga till språkkoden efter 
den vanliga URL-en. Som exempel hittar du den Italienska sidan under
*www.aros.org/it*, den Ryska på *www.aros.org/ru* och så vidare.

__ http://www.aros.org/fr/

AROS i nyheterna
----------------

Vi rekommenderar den här trevliga `recensionen`__ som Dmitar Butrovski har
skrivit på `OSnews.com`__. Det är utan tvekan en av de mest kompletta artiklar
som har skrivits om vårat fina operativsystem. Om du inte redan är bekant med
vad AROS är så får du antagligen en bra idé om det.

__ http://osnews.com/story.php?news_id=15819
__ http://osnews.com

Mjukvara
--------

Version 1.20 av den *VICE*, den berömda emulatorn av Commodores linje av
8-bitars datorer, finns nu tillgänglig för alla Amiga-plattformar inklusive AROS.
Du hittar den `här`__.

*WinAros* är en förinstallerad AROS-miljö installerad på en hårddisk-avbildning,
kompatibel med de välkända virtualiseringsmiljöerna QEMU och Microsoft
VirtualPC, båda fritt tillgängliga på Internet. Du kan ladda ner 
`QEMU Winaros här`__ och `QEMU VirtualPC här`__. Heinz-Raphael Reinke har också
skrivit en komplett guide över `AROS-installation på hårddisk`__ i PDF-format.
Den finns även på `Tyska`__ om du föredrar det. Du behöver Adobe Acrobat
Reader, FoxIt Reader eller aPDF/xPDF för att läsa dem.

*Installation Kit for AROS (IKAROS)* är en uppsättning med hårddisk-avbildningar
för olika virtualiseringsmiljöer, såsom QEMU och VMWare, redan partitionerade,
formatterade och färdiga att installera AROS på. Fördelarna med det är liten 
storlek på arkiven man laddar hem eftersom den inte behöver stora mängder med filer,
och möjligheten att installera nya, fräsha versioner av AROS. Det gör det enkelt
att testa nattliga kompileringar utan att behöva stöka med partitionering.
Instruktioner över hur man installerar medföljer.
Vänligen besök `Aros-Exec`__ för uppdateringar och nerladdning.

__ http://www.viceteam.org/amigaos.html
__ http://amidevcpp.amiga-world.de/WinAros/WinAros_Light_QEMU.zip
__ http://amidevcpp.amiga-world.de/WinAros/WinAros_Light_VPC.zip
__ http://amidevcpp.amiga-world.de/WinAros/Aros_HD_Install_English.pdf
__ http://amidevcpp.amiga-world.de/WinAros/Aros_HD_Installation.pdf
__ https://archives.aros-exec.org/?function=showfile&file=emulation/misc/arosik02.zip
