======
L�nkar
======

:Authors:   Aaron Digulla, Adam Chodorowski, Matthias Rustler 
:Copyright: Copyright � 1995-2007, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.


.. Contents::

AROS k�llor
===========

+ `Team AROS`__ 

  TeamAROS �r den ursprungliga supportgruppen f�r AROS.
  
+  `AROSWorld`__

  AROS Community hemsida, forum, nyheter, gallerier

+ `AROS software archive`__

+ `AROS Aminet Section`__

+ `AROS Polska`__

+ `AROS on ohloh.net`__

  Ohlow demonstrerar AROS-utvecklingens aktivitet p� ett snyggt grafiskt vis.

+ `Map of AROS users`__

+ `AROS for Amiga`__
  
  AfA OS byter ut AmigaOS core libraries med deras mer avancerade motsvarighet i AROS.
  
+ `AROS World`__
  En ny hemsida om AROS, avsedd f�r att vara en user community hemsida.

+ `AROS on WikiPedia`__

+ `AROS documentation on WikiBooks`__
  
__ http://www.teamaros.org/
__ https://www.arosworld.org/
__ http://archives.aros-exec.org/
__ http://aros.aminet.net/
__ http://www.aros.bbs.pl/
__ http://www.ohloh.net/projects/6056?p=AROS
__ http://www.frappr.com/arosusers
__ http://amidevcpp.amiga-world.de/afa_binarie_upload.php
__ http://arosworld.org
__ http://en.wikipedia.org/wiki/AROS_Research_Operating_System
__ http://en.wikibooks.org/wiki/Aros


Artiklar om AROS
================

===============================================  ==================  ==========
Titel                                            F�rfattare          Datum
===============================================  ==================  ==========
`"Onboard the Last Train to Amiga Neverland"`__  Dmitar Butrovski    2006-09-13
`"Test: AROS"`__ (in German mag. AmigaFuture)    Ingo Schmitz        2005-05-05
`"AROS"`__ (in German mag. Amiga-Magazin)        Martin Steigerwald  2003-09-13
`"If you like Amiga, you'll love AROS"`__        Elwood              Unknown   
`"AROS: Native AmigaOS For Your PC"`__           John Chandler       2001-10-21 
`"AROS: The Amiga Research Operating System`__   John Chandler       1999-10-02
===============================================  ==================  ==========

__ http://www.osnews.com/story.php?news_id=15819
__ http://www.amigafuture.de/kb.php?mode=article&k=1315&page_num=37&start=0
__ http://www.amiga-magazin.de/magazin/a09-03/aros/index.html
__ http://elwoodb.free.fr/articles/AROS/
__ http://www.suite101.com/article.cfm/amiga/82949 
__ http://www.suite101.com/article.cfm/amiga/26509

Om du k�nner till n�gon artikel om AROS som inte finns med, contact_ oss
s� vi kan l�gga till den. Tack.


Artiklar som n�mner AROS
========================

===============================================  ==============  ==========
Titel                                            F�rfattare      Datum
===============================================  ==============  ==========
`"Climbing the Kernel Mountain"`__               Emmanuel Marty  2002-08-13
`Interview with Martin Blom`__                   Johan Forsberg  Unknown
`"A Nudge In The Right Direction"`__             John Chandler   2002-07-02
`"What Are The Odds...?"`__                      John Chandler   2001-07-31
`"May Update"`__                                 John Chandler   2001-05-07
`"This Is Reality Control"`__                    John Chandler   2001-02-07
`"Open Amiga Foundation Update"`__               John Chandler   2000-07-02
`"Gui4Cli"`__                                    John Chandler   2000-03-01
`"And So It Begins..."`__                        John Chandler   2000-01-10
`"We're In This Together Now (Part II)"`__       John Chandler   1999-12-05
`"Open Source AmigaOS?"`__                       John Chandler   1999-03-01
===============================================  ==============  ==========

__ http://www.osnews.com/story.php?news_id=1532&page=1
__ http://www.kicker.nu/amigarulez/html/sections.php?op=viewarticle&artid=3
__ http://www.suite101.com/article.cfm/amiga/93270
__ http://www.suite101.com/article.cfm/amiga/76246
__ http://www.suite101.com/article.cfm/amiga/68505
__ http://www.suite101.com/article.cfm/amiga/59824
__ http://www.suite101.com/article.cfm/amiga/42265
__ http://www.suite101.com/article.cfm/amiga/34520
__ http://www.suite101.com/article.cfm/amiga/31482
__ http://www.suite101.com/article.cfm/amiga/29763
__ http://www.suite101.com/article.cfm/amiga/16364

Om du k�nner till n�gon artikel om AROS som inte finns med, contact_ oss
s� vi kan l�gga till den. Tack.

Utvecklarnas hemsidor
=====================

+ `Aaron Digulla`__
+ `Adam Chodorowski`__
+ `Henrik Berglund`__
+ `Johan Alfredsson`__
+ `Lennard voor den Dag`__
+ `Martin Steigerwald`__
+ `Matt 'Crazy' Parsons`__
+ `Matthias Rustler`__
+ `Michal Schulz`__
+ `Nic Andrews`__
+ `Oliver Brunner`__
+ `Olivier Adam`__
+ `Robert Norris`__
+ `Sebastian Rittau`__


__ http://www.philmann-dark.de/
__ http://www.chodorowski.com/
__ http://www.mds.mdh.se/~adb94hbd/
__ http://www.dtek.chalmers.se/~d95duvan/
__ http://www.xs4all.nl/~ldp/
__ http://www.lichtvoll.de
__ http://www.troubled-mind.com
__ http://www.mazze-online.de/
__ http://msaros.blogspot.com
__ http://kalamatee.blogspot.com/
__ http://homes.hallertau.net/~oli/
__ http://reziztanzia.free.fr/
__ http://cataclysm.cx/
__ http://www.in-berlin.de/User/jroger/index.html


�vrigt
======

+ `Back to the Roots`__

  .. Image:: ./images/bttr.jpeg

  En suver�n nostalgi-sida d�r du kan hitta licensierade och fria Amiga-spel.


__ http://www.back2roots.org/


.. _contact: contact
