==================
Kontaktinformation
==================

:Authors:   Adam Chodorowski, Matthias Rustler 
:Copyright: Copyright © 1995-2009, The AROS Development Team
:Version:   $Revision$
:Date:      $Date$
:Status:    Done.

.. Contents::


Kontakperson
============
Den primära kontaktpersonen för teamet som utvecklar AROS är Aaron "Optimizer"
Digulla. Om du vill ha kontakt med AROS som projekt, till exempel för att diskutera
sponsoravtal eller andra former av samarbete, så är det personen att kontakta.
Du kan nå honom genom att skicka email till `digulla@aros.org`__.

__ mailto:digulla@aros.org


Mailinglistor
=============

Det finns ett antal AROS-relaterade mailinglistor, vilka är de viktigaste kanalerna
för information och diskussion om AROS för utvecklare. Följande mailinglistor finns
tillgängliga:

+ `AROS Developer`__

  Det här är listan för utvecklare där diskussioner om utvecklingen av AROS sker.
  Här postas också statusen från den nattliga kompileringen av AROS. Det är 
  **starkt** rekommenderat att utvecklare går med i den här listan eftersom det
  annars är svårt att hålla sig uppdaterad med den senaste utvecklingen.
  Eftersom det inte finns så många utvecklare inom AROS, så är mängden email
  ganska liten men den kan bli ganska hög om en het diskussion kommer igång.

  .. Note:: Begäran om prenumeration på den här listan hanteras inte automatiskt
            utan varje begäran kontrolleras av listans administratörer. Detta
            innebär att det kan ta ett litet tag från det att du skickar in 
            en begäran tills dess att du blir en medlem.
  
+ `AROS CVS`__

  På denna lista för utvecklare postas loggar från Subversion-servern så fort något
  sänder in ändringar ("commit"). I motsats till den dagliga samlings-loggen som 
  postas på AROS Developer-listan, där varje mail innehåller hela dagens aktiviteter
  på Subversion-servern, så skickas det separata email för varje insänd ändring
  *omedelbart* för varje loggad aktivitet. Så om du vill ha nästan realtids-information
  om vad som händer på Subversion-servern så är det här listan för dig.
  Volymen av mail på denna lista kan vara ganska hög.

+ `AROS Website`__

  Skriptsystemet som skapar hemsidan skickar mail till den här listan.
  De som jobbar med dokumentationen eller kan laga saker om  något händer
  med websidan bör prenumerera på denna.

Följ länkarna till de administrativa sidorna för information om hur man
prenumererar, avbryter prenumerationerer, listarkiv och andra användbara
funktioner.

__ https://mail.aros.org/mailman/listinfo/aros-dev
__ http://lists.sourceforge.net/mailman/listinfo/aros-cvs
__ http://lists.sourceforge.net/mailman/listinfo/aros-website

.. _`buggdatabasen`: http://sourceforge.net/tracker/?atid=439463&group_id=43586&func=browse


Forum
=====

AROS-Exec__ är den officella community-portalen för AROS. Här finner du de
senaste nyheterna om AROS, diskussionsforum, bildgallerier och mycket mer. Det
är den perfekta mötesplatsen för AROS-användare från hela världen.

__ https://www.arosworld.org/

IRC-Kanaler
===========

Det finns en officiell IRC-kanal för AROS, föga förvånande döpt till `#aros`__, på
FreeNode__-nätverket. Vänligen anslut till `irc.freenode.net`__ som vidarebefodrar 
dig till en server nära dig. Den är till för att diskutera allt möjligt som är relaterat
med AROS inklusive utveckling och planer att ta över världen. Vid sällsynta tillfällen
när det är väldigt mycket prat i huvudkanalen flyttar diskussioner relaterade till
utveckling till `#aros.dev`__.

__ irc://irc.freenode.net/aros
__ http://www.freenode.net/
__ irc://irc.freenode.net/
__ irc://irc.freenode.net/aros.dev
